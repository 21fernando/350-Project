module IO(
    input clk,
    input [31:0] IO_read_1,
    input [31:0] IO_read_2,
    input [31:0] IO_read_3,
    input [31:0] IO_read_4,
    input [31:0] IO_read_5,
    output [31:0] IO_write_1,
    output [31:0] IO_write_2,
    output [31:0] IO_write_3,
    output [31:0] IO_write_4,
    output [31:0] IO_write_5,
    output [4:0] IO_wEn);

    

endmodule